package Constants;
    
    //Screen size
    parameter SCREEN_HEIGHT = 9'd480;
    parameter SCREEN_WIDTH = 10'd640;

    //Obstacle sizes
    parameter OBSTACLE_MIN_Y = 6'd50;
    parameter OBSTACLE_MAX_Y = 8'd200;
    parameter OBSTACLE_MAX_DISTANCE = 10'd680;
    parameter OBSTACLE_WIDTH = 6'd40;
    parameter TIME_TO_OBSTACLE = 6'd50; //tbd

    //Bird Width
    
    parameter BIRD_WIDTH = 6'40; 
